
`define	ADDI			3'b001
`define	ADD			3'b010
`define	BNE			3'b011
`define	BEQ			3'b100
`define	LDI			3'b101
`define	MUL			3'b110