
`define	RA			3'b101
`define	RADDI			3'b001
`define	RADD			3'b010	
`define	RSUBI			6'b011
`define	RSUB			6'b100				
`define	RMUL			3'b110
